-- [B: 30|PDF: 38] Chapter 1 "Fundamental Concepts" - Ex. 8
-- Task: 

-- Answer:
