-- [B: 30|PDF: 38] Chapter 1 "Fundamental Concepts" - Ex. 4
-- Task: 
-- 4. [➊ 1.5] Rewrite the following decimal literals as hexadecimal literals.

-- Answer:
-- 0000 0000 0000 0000
--                | |1
--                | 16
--                |256
--                4096

-- Decimal  -> HEX
-- 1        -> x0001  x1
-- 34       -> x0022
-- 256.0    -> x0100.0000
-- 0.5      -> x0000.8  x0000.8000  16x0000.8
