-- [B: 94|PDF:102] Chapter 3 "Sequential Statements" - Ex. 1
-- Task: 

-- Answer: