-- [B:135|PDF:143] Chapter 4 "Composite Data Types and Operations" - Ex. 1
-- Task: 

-- Answer:
