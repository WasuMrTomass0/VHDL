-- [B:243|PDF:251] Chapter 6 "Subprograms" - Ex. 8
-- Task: 

-- Answer:
