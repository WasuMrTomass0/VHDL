-- [B: 30|PDF: 38] Chapter 1 "Fundamental Concepts" - Ex. 4
-- Task: 

-- Answer: