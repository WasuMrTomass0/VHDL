-- [B:205|PDF:213] Chapter 5 "Basic Modeling Constructs" - Ex. 15
-- Task: 

-- Answer:
